module sbox_32bit
(									
    input	[31:0]	a_i,
    output	logic[31:0]	d_o
);

	sbox_8bit s0(a_i[7:0],   d_o[7:0]);
	sbox_8bit s1(a_i[15:8],  d_o[15:8]);
	sbox_8bit s2(a_i[23:16], d_o[23:16]);
	sbox_8bit s3(a_i[31:24], d_o[31:24]);
	
endmodule

module sbox_8bit
(										
    input	[7:0]	a_i,
    output	logic[7:0]	d_o
);
always_comb
	case(a_i)
		8'h00:	d_o	=	8'hd6;
		8'h01:	d_o	=	8'h90;
		8'h02:	d_o	=	8'he9;
		8'h03:	d_o	=	8'hfe;
		8'h04:	d_o	=	8'hcc;
		8'h05:	d_o	=	8'he1;
		8'h06:	d_o	=	8'h3d;
		8'h07:	d_o	=	8'hb7;
		8'h08:	d_o	=	8'h16;
		8'h09:	d_o	=	8'hb6;
		8'h0a:	d_o	=	8'h14;
		8'h0b:	d_o	=	8'hc2;
		8'h0c:	d_o	=	8'h28;
		8'h0d:	d_o	=	8'hfb;
		8'h0e:	d_o	=	8'h2c;
		8'h0f:	d_o	=	8'h05;
		8'h10:	d_o	=	8'h2b;
		8'h11:	d_o	=	8'h67;
		8'h12:	d_o	=	8'h9a;
		8'h13:	d_o	=	8'h76;
		8'h14:	d_o	=	8'h2a;
		8'h15:	d_o	=	8'hbe;
		8'h16:	d_o	=	8'h04;
		8'h17:	d_o	=	8'hc3;
		8'h18:	d_o	=	8'haa;
		8'h19:	d_o	=	8'h44;
		8'h1a:	d_o	=	8'h13;
		8'h1b:	d_o	=	8'h26;
		8'h1c:	d_o	=	8'h49;
		8'h1d:	d_o	=	8'h86;
		8'h1e:	d_o	=	8'h06;
		8'h1f:	d_o	=	8'h99;
		8'h20:	d_o	=	8'h9c;
		8'h21:	d_o	=	8'h42;
		8'h22:	d_o	=	8'h50;
		8'h23:	d_o	=	8'hf4;
		8'h24:	d_o	=	8'h91;
		8'h25:	d_o	=	8'hef;
		8'h26:	d_o	=	8'h98;
		8'h27:	d_o	=	8'h7a;
		8'h28:	d_o	=	8'h33;
		8'h29:	d_o	=	8'h54;
		8'h2a:	d_o	=	8'h0b;
		8'h2b:	d_o	=	8'h43;
		8'h2c:	d_o	=	8'hed;
		8'h2d:	d_o	=	8'hcf;
		8'h2e:	d_o	=	8'hac;
		8'h2f:	d_o	=	8'h62;
		8'h30:	d_o	=	8'he4;
		8'h31:	d_o	=	8'hb3;
		8'h32:	d_o	=	8'h1c;
		8'h33:	d_o	=	8'ha9;
		8'h34:	d_o	=	8'hc9;
		8'h35:	d_o	=	8'h08;
		8'h36:	d_o	=	8'he8;
		8'h37:	d_o	=	8'h95;
		8'h38:	d_o	=	8'h80;
		8'h39:	d_o	=	8'hdf;
		8'h3a:	d_o	=	8'h94;
		8'h3b:	d_o	=	8'hfa;
		8'h3c:	d_o	=	8'h75;
		8'h3d:	d_o	=	8'h8f;
		8'h3e:	d_o	=	8'h3f;
		8'h3f:	d_o	=	8'ha6;
		8'h40:	d_o	=	8'h47;
		8'h41:	d_o	=	8'h07;
		8'h42:	d_o	=	8'ha7;
		8'h43:	d_o	=	8'hfc;
		8'h44:	d_o	=	8'hf3;
		8'h45:	d_o	=	8'h73;
		8'h46:	d_o	=	8'h17;
		8'h47:	d_o	=	8'hba;
		8'h48:	d_o	=	8'h83;
		8'h49:	d_o	=	8'h59;
		8'h4a:	d_o	=	8'h3c;
		8'h4b:	d_o	=	8'h19;
		8'h4c:	d_o	=	8'he6;
		8'h4d:	d_o	=	8'h85;
		8'h4e:	d_o	=	8'h4f;
		8'h4f:	d_o	=	8'ha8;
		8'h50:	d_o	=	8'h68;
		8'h51:	d_o	=	8'h6b;
		8'h52:	d_o	=	8'h81;
		8'h53:	d_o	=	8'hb2;
		8'h54:	d_o	=	8'h71;
		8'h55:	d_o	=	8'h64;
		8'h56:	d_o	=	8'hda;
		8'h57:	d_o	=	8'h8b;
		8'h58:	d_o	=	8'hf8;
		8'h59:	d_o	=	8'heb;
		8'h5a:	d_o	=	8'h0f;
		8'h5b:	d_o	=	8'h4b;
		8'h5c:	d_o	=	8'h70;
		8'h5d:	d_o	=	8'h56;
		8'h5e:	d_o	=	8'h9d;
		8'h5f:	d_o	=	8'h35;
		8'h60:	d_o	=	8'h1e;
		8'h61:	d_o	=	8'h24;
		8'h62:	d_o	=	8'h0e;
		8'h63:	d_o	=	8'h5e;
		8'h64:	d_o	=	8'h63;
		8'h65:	d_o	=	8'h58;
		8'h66:	d_o	=	8'hd1;
		8'h67:	d_o	=	8'ha2;
		8'h68:	d_o	=	8'h25;
		8'h69:	d_o	=	8'h22;
		8'h6a:	d_o	=	8'h7c;
		8'h6b:	d_o	=	8'h3b;
		8'h6c:	d_o	=	8'h01;
		8'h6d:	d_o	=	8'h21;
		8'h6e:	d_o	=	8'h78;
		8'h6f:	d_o	=	8'h87;
		8'h70:	d_o	=	8'hd4;
		8'h71:	d_o	=	8'h00;
		8'h72:	d_o	=	8'h46;
		8'h73:	d_o	=	8'h57;
		8'h74:	d_o	=	8'h9f;
		8'h75:	d_o	=	8'hd3;
		8'h76:	d_o	=	8'h27;
		8'h77:	d_o	=	8'h52;
		8'h78:	d_o	=	8'h4c;
		8'h79:	d_o	=	8'h36;
		8'h7a:	d_o	=	8'h02;
		8'h7b:	d_o	=	8'he7;
		8'h7c:	d_o	=	8'ha0;
		8'h7d:	d_o	=	8'hc4;
		8'h7e:	d_o	=	8'hc8;
		8'h7f:	d_o	=	8'h9e;
		8'h80:	d_o	=	8'hea;
		8'h81:	d_o	=	8'hbf;
		8'h82:	d_o	=	8'h8a;
		8'h83:	d_o	=	8'hd2;
		8'h84:	d_o	=	8'h40;
		8'h85:	d_o	=	8'hc7;
		8'h86:	d_o	=	8'h38;
		8'h87:	d_o	=	8'hb5;
		8'h88:	d_o	=	8'ha3;
		8'h89:	d_o	=	8'hf7;
		8'h8a:	d_o	=	8'hf2;
		8'h8b:	d_o	=	8'hce;
		8'h8c:	d_o	=	8'hf9;
		8'h8d:	d_o	=	8'h61;
		8'h8e:	d_o	=	8'h15;
		8'h8f:	d_o	=	8'ha1;
		8'h90:	d_o	=	8'he0;
		8'h91:	d_o	=	8'hae;
		8'h92:	d_o	=	8'h5d;
		8'h93:	d_o	=	8'ha4;
		8'h94:	d_o	=	8'h9b;
		8'h95:	d_o	=	8'h34;
		8'h96:	d_o	=	8'h1a;
		8'h97:	d_o	=	8'h55;
		8'h98:	d_o	=	8'had;
		8'h99:	d_o	=	8'h93;
		8'h9a:	d_o	=	8'h32;
		8'h9b:	d_o	=	8'h30;
		8'h9c:	d_o	=	8'hf5;
		8'h9d:	d_o	=	8'h8c;
		8'h9e:	d_o	=	8'hb1;
		8'h9f:	d_o	=	8'he3;
		8'ha0:	d_o	=	8'h1d;
		8'ha1:	d_o	=	8'hf6;
		8'ha2:	d_o	=	8'he2;
		8'ha3:	d_o	=	8'h2e;
		8'ha4:	d_o	=	8'h82;
		8'ha5:	d_o	=	8'h66;
		8'ha6:	d_o	=	8'hca;
		8'ha7:	d_o	=	8'h60;
		8'ha8:	d_o	=	8'hc0;
		8'ha9:	d_o	=	8'h29;
		8'haa:	d_o	=	8'h23;
		8'hab:	d_o	=	8'hab;
		8'hac:	d_o	=	8'h0d;
		8'had:	d_o	=	8'h53;
		8'hae:	d_o	=	8'h4e;
		8'haf:	d_o	=	8'h6f;
		8'hb0:	d_o	=	8'hd5;
		8'hb1:	d_o	=	8'hdb;
		8'hb2:	d_o	=	8'h37;
		8'hb3:	d_o	=	8'h45;
		8'hb4:	d_o	=	8'hde;
		8'hb5:	d_o	=	8'hfd;
		8'hb6:	d_o	=	8'h8e;
		8'hb7:	d_o	=	8'h2f;
		8'hb8:	d_o	=	8'h03;
		8'hb9:	d_o	=	8'hff;
		8'hba:	d_o	=	8'h6a;
		8'hbb:	d_o	=	8'h72;
		8'hbc:	d_o	=	8'h6d;
		8'hbd:	d_o	=	8'h6c;
		8'hbe:	d_o	=	8'h5b;
		8'hbf:	d_o	=	8'h51;
		8'hc0:	d_o	=	8'h8d;
		8'hc1:	d_o	=	8'h1b;
		8'hc2:	d_o	=	8'haf;
		8'hc3:	d_o	=	8'h92;
		8'hc4:	d_o	=	8'hbb;
		8'hc5:	d_o	=	8'hdd;
		8'hc6:	d_o	=	8'hbc;
		8'hc7:	d_o	=	8'h7f;
		8'hc8:	d_o	=	8'h11;
		8'hc9:	d_o	=	8'hd9;
		8'hca:	d_o	=	8'h5c;
		8'hcb:	d_o	=	8'h41;
		8'hcc:	d_o	=	8'h1f;
		8'hcd:	d_o	=	8'h10;
		8'hce:	d_o	=	8'h5a;
		8'hcf:	d_o	=	8'hd8;
		8'hd0:	d_o	=	8'h0a;
		8'hd1:	d_o	=	8'hc1;
		8'hd2:	d_o	=	8'h31;
		8'hd3:	d_o	=	8'h88;
		8'hd4:	d_o	=	8'ha5;
		8'hd5:	d_o	=	8'hcd;
		8'hd6:	d_o	=	8'h7b;
		8'hd7:	d_o	=	8'hbd;
		8'hd8:	d_o	=	8'h2d;
		8'hd9:	d_o	=	8'h74;
		8'hda:	d_o	=	8'hd0;
		8'hdb:	d_o	=	8'h12;
		8'hdc:	d_o	=	8'hb8;
		8'hdd:	d_o	=	8'he5;
		8'hde:	d_o	=	8'hb4;
		8'hdf:	d_o	=	8'hb0;
		8'he0:	d_o	=	8'h89;
		8'he1:	d_o	=	8'h69;
		8'he2:	d_o	=	8'h97;
		8'he3:	d_o	=	8'h4a;
		8'he4:	d_o	=	8'h0c;
		8'he5:	d_o	=	8'h96;
		8'he6:	d_o	=	8'h77;
		8'he7:	d_o	=	8'h7e;
		8'he8:	d_o	=	8'h65;
		8'he9:	d_o	=	8'hb9;
		8'hea:	d_o	=	8'hf1;
		8'heb:	d_o	=	8'h09;
		8'hec:	d_o	=	8'hc5;
		8'hed:	d_o	=	8'h6e;
		8'hee:	d_o	=	8'hc6;
		8'hef:	d_o	=	8'h84;
		8'hf0:	d_o	=	8'h18;
		8'hf1:	d_o	=	8'hf0;
		8'hf2:	d_o	=	8'h7d;
		8'hf3:	d_o	=	8'hec;
		8'hf4:	d_o	=	8'h3a;
		8'hf5:	d_o	=	8'hdc;
		8'hf6:	d_o	=	8'h4d;
		8'hf7:	d_o	=	8'h20;
		8'hf8:	d_o	=	8'h79;
		8'hf9:	d_o	=	8'hee;
		8'hfa:	d_o	=	8'h5f;
		8'hfb:	d_o	=	8'h3e;
		8'hfc:	d_o	=	8'hd7;
		8'hfd:	d_o	=	8'hcb;
		8'hfe:	d_o	=	8'h39;
		8'hff:	d_o	=	8'h48;
	endcase
endmodule